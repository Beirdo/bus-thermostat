SPWM2 (PSpice format)
**************************************
**  This file was created by TINA   **
**         www.tina.com             ** 
**      (c) DesignSoft, Inc.        **          
**     www.designsoftware.com       **
**************************************
.LIB "C:\Program Files (x86)\DesignSoft\Tina 9 - TI\EXAMPLES\SPICE\TSPICE.LIB"
.LIB "C:\Program Files (x86)\DesignSoft\Tina 9 - TI\SPICELIB\Operational Amplifiers.LIB"
.LIB
.TEMP 27
.AC DEC 20 10 1MEG
.TRAN 400U 200M UIC

.OPTIONS ABSTOL=1P ITL1=150 ITL2=20 ITL4=10 TRTOL=7 
.PROBE V([VF6]) V([VF4]) V([VF1]) V([VF3]) V([VF5])
.PROBE V([VF2])

V8          4 0 12
V1          21 0 12
V3          0 26 6
V2          20 0 6
V7          0 33 6
V6          14 0 6
V4          0 38 6
V5          37 0 6
LM1_1       1 2 437U
LM1_2       VF6 0 874U
KM1         LM1_1       LM1_2       1.4142135624
L1          6 VF4 1.5M IC=0 
XU15        8 VF1 IC_7417_0
XU14        10 VF3 IC_7417_0
R18         11 12 10K 
R17         11 13 10K 
XU13        0 11 14 0 13 LMV651_0
XU12        15 10 14 0 10 LMV651_0
XU11        16 13 14 0 15 LMV651_0
R23         17 VF2 10K 
R22         17 16 10K 
XU10        0 17 14 0 16 LMV651_0
XU7         19 8 20 0 8 LMV651_0
R16         21 22 100MEG 
R11         23 0 10K 
XP2          24 23 VF5  PotMeter PARAMS: Res=50K Percent=10M
XU5         22 23 20 26 VF5 LMV651_0
R5          22 0 1.2MEG 
C3          27 22 10P IC=0 
XU4         28 27 21 0 27 LMV651_0
XU1          28 29 28   21   30   31   21   0  CA555 ; Timer
C1          28 0 100P 
C2          29 0 10N 
R1          28 31 143K 
R2          21 31 1K 
XU9         VF2 12 20 0 19 LMV651_0
XU8         VF5 12 20 26 12 LMV651_0
R15         32 0 10K 
R3          32 VF2 220K 
XU6         34 32 14 33 VF2 LMV651_0
XU2         0 35 37 38 36 LMV651_0
R14         35 34 10K 
R6          36 35 560K 
C5          0 34 2.2U IC=0 
R9          39 34 1.21K 
C4          0 39 2.2U IC=0 
R4          40 39 1.21K 
C6          0 40 2.2U IC=0 
R13         36 40 1.21K 
R12         VF6 6 10 
C13         0 VF4 68U IC=0 
R10         41 1 200 
C11         41 4 10U IC=0 
C10         0 41 10U IC=0 
R7          42 43 200 
R8          44 45 200 
MT2         2 45 0 0  ME_IRF540_N_1 NRD=0 NRS=0 
MT1         4 43 2 2  ME_IRF540_N_1 NRD=0 NRS=0 
C9          4 0 100N IC=0 
C8          46 2 100N IC=0 
XU3         2 VF1 42 46 VF3 44 4 0 UCC27211_TRANS

.MODEL ME_IRF540_N_1 NMOS( LEVEL=3 VTO=3.134 KP=20.59U PHI=600M GAMMA=0 TOX=100N 
+      UO=600 VMAX=0 DELTA=0 THETA=0 ETA=0 
+      L=2U W=940M RD=22.52M RS=21.34M RG=5.557 
+      RB=0 RDS=444.4K IS=2.848P N=1 PB=800M 
+      CBD=2.422N CBS=0 MJ=500M TT=142N CGSO=1.144N 
+      CGDO=443.8P CGBO=0 KF=0 AF=1 )

.LIB "C:\Program Files (x86)\DesignSoft\Tina 9 - TI\SPICELIB\NSC.LIB"
* END MODEL LMV641

* BEGIN MODEL LMV651
*//////////////////////////////////////////////////////////////////////
* (C) NATIONAL SEMICONDUCTOR, CORPORATION.
* MODELS DEVELOPED AND UNDER COPYRIGHT BY:
* NATIONAL SEMICONDUCTOR, CORPORATION.
*/////////////////////////////////////////////////////////////////////
* LEGAL NOTICE:
* THE MODEL MAY BE COPIED, AND DISTRIBUTED WITHOUT ANY MODIFICATIONS;
* HOWEVER, RESELLING OR LICENSING THE MATERIAL IS ILLEGAL.
* WE RESERVE THE RIGHT TO MAKE CHANGES TO THE MODEL WITHOUT PRIOR NOTICE.
* PSPICE MODELS ARE PROVIDED "AS IS, WITH NO WARRANTY OF ANY KIND"
*////////////////////////////////////////////////////////////////////
* MODEL FEATURES INCLUDE OUTPUT SWING, OUTPUT CURRENT THRU
* THE SUPPLY RAILS, OUTPUT SWING VS IO, OUTPUT CURRENT LIMIT,
* OPEN LOOP GAIN AND PHASE, SLEW RATE, COMMON MODE REJECTION
* WITH FREQ EFFECTS, POWER SUPPLY REJECTION WITH FREQ EFFECTS,
* INPUT VOLTAGE NOISE WITH 1/F, INPUT CURRENT NOISE, INPUT
* CAPACITANCE, INPUT BIAS CURRENT, INPUT COMMON MODE RANGE,
* INPUT OFFSET, HIGH CLOAD EFFECTS, AND QUIESCENT CURRENT
* VS VOLTAGE AND TEMPERATURE.
*///////////////////////////////////////////////////////////////
* MODEL TEMP RANGE IS -40 TO +125 DEG C.
* NOTE THAT MODEL IS FUNCTIONAL OVER THIS RANGE BUT NOT ALL
* PARAMETERS TRACK THOSE OF THE REAL PART.
*////////////////////////////////////////////////////////////
* PINOUT ORDER +IN -IN V+ V- OUT
* PINOUT ORDER  1   3   5  2  4
.SUBCKT LMV651_0  1 3 5 2 4
Q12 6 7 8 QP
Q13 9 9 10 QP
Q14 11 11 9 QP
Q15 8 12 10 QP
Q17 13 8 14 QOP
Q18 15 15 16 QN
Q19 16 16 17 QN
Q20 6 18 19 QN
Q21 20 6 21 QON
Q22 8 15 6 QN
R10 18 22 100
R11 12 23 100
R12 14 5 50
R13 2 21 4
G1 6 19 24 25 -2E-4
R16 24 26 100
C2 26 4 17E-12
R17 7 11 50
R18 19 17 4
D5 4 5 DD
D6 2 4 DD
E2 19 0 2 0 1
E3 10 0 5 0 1
I12 5 2 105E-6
G4 24 25 27 28 2E-3
R40 24 25 9E5
E14 25 19 10 19 0.5
D11 24 10 DD
D12 19 24 DD
R41 20 4 2
R42 4 13 4
Q23 8 29 10 QP
Q24 15 30 10 QP
Q25 6 31 19 QN
Q26 7 32 19 QN
Q33 33 34 10 QP
R45 35 36 1
R46 37 36 1
R47 38 39 7E3
R49 19 27 425
R50 19 28 425
R51 40 41 7E3
Q35 41 41 42 QP
Q37 42 42 41 QN
D13 42 10 DD
D14 41 10 DD
D15 43 42 DD
D16 43 41 DD
V10 39 42 -0.07E-3
D17 44 0 DIN
D18 45 0 DIN
I14 0 44 0.1E-3
I15 0 45 0.1E-3
C13 38 0 3E-12
C14 3 0 3E-12
D19 46 0 DVN
D20 47 0 DVN
I16 0 46 0.1E-3
I17 0 47 0.1E-3
E15 40 3 46 47 1.75
G5 38 40 44 45 3.6E-5
E16 49 0 10 0 1
E17 50 0 19 0 1
E18 51 0 52 0 1
R56 49 53 1E6
R57 50 54 1E6
R58 51 55 1E6
R59 0 53 100
R60 0 54 100
R61 0 55 100
E19 56 1 55 0 -47E-3
R62 57 52 1E3
R63 52 58 1E3
C15 49 53 1E-12
C16 50 54 1E-12
C17 51 55 70E-12
E20 59 56 54 0 0.25
E21 38 59 53 0 -0.20
C19 27 28 8E-12
G6 34 10 60 0 0.68E-6
G7 29 10 60 0 3.4E-7
G8 30 10 60 0 1.45E-7
G9 19 31 60 0 1.7E-7
G10 19 32 60 0 7.25E-8
R64 0 60 1E12
R132 4 24 1E8
I18 38 0 80E-9
I19 3 0 80E-9
V53 43 19 0.07
V54 33 36 0.1
G12 38 40 61 0 8E-6
R136 0 61 12E3
R137 0 61 12E3
R138 1 56 1E9
R139 56 59 1E9
R140 59 38 1E9
E54 58 0 38 0 1
E55 57 0 40 0 1
C23 38 40 0.25E-12
E72 22 19 21 2 3.5
E73 23 10 14 10 0.75
M61 28 42 35 35 MIP L=2U W=150U
M62 27 41 37 37 MIP L=2U W=150U
V55 60 0 1
R141 2 5 1E6
G13 5 2 62 0 -2E-4
I20 0 63 1E-3
D21 63 0 DD
V56 63 62 0.65
R143 0 62 1E6
.MODEL QON NPN VAF=40
.MODEL QOP PNP VAF=40
.MODEL MIP PMOS KP=600U VTO=-0.7
.MODEL DD D
.MODEL QN NPN
.MODEL QP PNP
.MODEL DVN D KF=0.7E-16
.MODEL DIN D KF=8E-17
.ENDS


.LIB "C:\Program Files (x86)\DesignSoft\Tina 9 - TI\SPICELIB\UCC27211_TRANS.LIB"
* SUBCKT: UCC27211_TRANS encrypted macro, content not displayed


.SUBCKT IC_7417_0 1A 1B
UNoname     BUF $G_DPWR $G_DGND  1A 1B  U_SN7407_1 IO_STD_OC
.MODEL U_SN7407_1 UGATE( TPLHTY=10N TPHLTY=10N )
.ENDS


.END
